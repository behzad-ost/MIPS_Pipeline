library verilog;
use verilog.vl_types.all;
entity test_CPU is
end test_CPU;
